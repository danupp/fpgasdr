// clkctrl_main.v

// Generated using ACDS version 15.1 193

`timescale 1 ps / 1 ps
module clkctrl_main (
		input  wire  inclk1x,   //  altclkctrl_input.inclk1x
		input  wire  inclk0x,   //                  .inclk0x
		input  wire  clkselect, //                  .clkselect
		output wire  outclk     // altclkctrl_output.outclk
	);

	clkctrl_main_altclkctrl_0 altclkctrl_0 (
		.inclk1x   (inclk1x),   //  altclkctrl_input.inclk1x
		.inclk0x   (inclk0x),   //                  .inclk0x
		.clkselect (clkselect), //                  .clkselect
		.outclk    (outclk)     // altclkctrl_output.outclk
	);

endmodule
