library ieee;
use ieee.std_logic_1164.ALL;
use ieee.std_logic_unsigned.ALL;
use ieee.numeric_std.ALL;

entity down_dec is
	port (Data_in : in std_logic_vector(23 downto 0);
			Data_out_I : out std_logic_vector(23 downto 0);
			Data_out_Q : out std_logic_vector(23 downto 0);
			clk_in : in std_logic; 
			clk_sample : in std_logic; 
			rx_att : in std_logic_vector(1 downto 0);
			clk_out : out std_logic
			);
end down_dec;

architecture down_dec_arch of down_dec is
	
type longbuffer is array (0 to 257) of signed (23 downto 0);
type filt_type is array (0 to 247) of signed (23 downto 0);

signal Ia : longbuffer;
signal Qa : longbuffer;

constant filtkoeff : filt_type :=

-- Scilab:
-->[v,a,f] = wfir ('lp', 496, [12/1250 0], 'hn', 20);
--> round(v*2^28)

	("000000000000000000000000",
    "000000000000000000001010",
    "000000000000000000101100",
    "000000000000000001101000",
    "000000000000000011000001",
    "000000000000000100111001",
    "000000000000000111010010",
    "000000000000001010001101",
    "000000000000001101101011",
    "000000000000010001101100",
    "000000000000010110001110",
    "000000000000011011010000",
    "000000000000100000110000",
    "000000000000100110101011",
    "000000000000101100111101",
    "000000000000110011100011",
    "000000000000111010011000",
    "000000000001000001010110",
    "000000000001001000010110",
    "000000000001001111010011",
    "000000000001010110000101",
    "000000000001011100100100",
    "000000000001100010101001",
    "000000000001101000001010",
    "000000000001101100111111",
    "000000000001110000111111",
    "000000000001110100000001",
    "000000000001110101111011",
    "000000000001110110100100",
    "000000000001110101110010",
    "000000000001110011011101",
    "000000000001101111011100",
    "000000000001101001100110",
    "000000000001100001110010",
    "000000000001010111111010",
    "000000000001001011110110",
    "000000000000111101011111",
    "000000000000101100110000",
    "000000000000011001100100",
    "000000000000000011110111",
    "111111111111101011100111",
    "111111111111010000110001",
    "111111111110110011010101",
    "111111111110010011010100",
    "111111111101110000101111",
    "111111111101001011101001",
    "111111111100100100001000",
    "111111111011111010010000",
    "111111111011001110001010",
    "111111111010011111111111",
    "111111111001101111111000",
    "111111111000111110000001",
    "111111111000001010101001",
    "111111110111010101111101",
    "111111110110100000001110",
    "111111110101101001101101",
    "111111110100110010101110",
    "111111110011111011100100",
    "111111110011000100100101",
    "111111110010001110001000",
    "111111110001011000100100",
    "111111110000100100010011",
    "111111101111110001101101",
    "111111101111000001001101",
    "111111101110010011001101",
    "111111101101101000001010",
    "111111101101000000011110",
    "111111101100011100100111",
    "111111101011111100111111",
    "111111101011100010000010",
    "111111101011001100001101",
    "111111101010111011111011",
    "111111101010110001100101",
    "111111101010101101100110",
    "111111101010110000010110",
    "111111101010111010001100",
    "111111101011001011100000",
    "111111101011100100100110",
    "111111101100000101110000",
    "111111101100101111010000",
    "111111101101100001010101",
    "111111101110011100001011",
    "111111101111011111111101",
    "111111110000101100110011",
    "111111110010000010110010",
    "111111110011100001111101",
    "111111110101001010010010",
    "111111110110111011101110",
    "111111111000110110001010",
    "111111111010111001011100",
    "111111111101000101010111",
    "111111111111011001101010",
    "000000000001110110000000",
    "000000000100011010000010",
    "000000000111000101010011",
    "000000001001110111010110",
    "000000001100101111101001",
    "000000001111101101100100",
    "000000010010110000011111",
    "000000010101110111101110",
    "000000011001000010100000",
    "000000011100010000000011",
    "000000011111011111100001",
    "000000100010110000000001",
    "000000100110000000101000",
    "000000101001010000011000",
    "000000101100011110010000",
    "000000101111101001001111",
    "000000110010110000010000",
    "000000110101110010001101",
    "000000111000101110000001",
    "000000111011100010100010",
    "000000111110001110100111",
    "000001000000110001001001",
    "000001000011001000111101",
    "000001000101010100111011",
    "000001000111010011111011",
    "000001001001000100110100",
    "000001001010100110100010",
    "000001001011110111111110",
    "000001001100111000001000",
    "000001001101100101111111",
    "000001001110000000100110",
    "000001001110000111000011",
    "000001001101111000011111",
    "000001001101010100001000",
    "000001001100011001001111",
    "000001001011000111001011",
    "000001001001011101010111",
    "000001000111011011010010",
    "000001000101000000100011",
    "000001000010001100110110",
    "000000111110111111111100",
    "000000111011011001101111",
    "000000110111011010001100",
    "000000110011000001011011",
    "000000101110001111100111",
    "000000101001000101000101",
    "000000100011100010010001",
    "000000011101100111101111",
    "000000010111010110001000",
    "000000010000101110010001",
    "000000001001110001000011",
    "000000000010011111100000",
    "111111111010111010110011",
    "111111110011000100001101",
    "111111101010111101001001",
    "111111100010100111000110",
    "111111011010000011101101",
    "111111010001010100101111",
    "111111001000011100000001",
    "111110111111011011100001",
    "111110110110010101010010",
    "111110101101001011100000",
    "111110100100000000011001",
    "111110011010110110010100",
    "111110010001101111101011",
    "111110001000101110111101",
    "111101111111110110101101",
    "111101110111001001100010",
    "111101101110101010001000",
    "111101100110011011001011",
    "111101011110011111011010",
    "111101010110111001100111",
    "111101001111101100100011",
    "111101001000111011000000",
    "111101000010100111110001",
    "111100111100110101100111",
    "111100110111100111010001",
    "111100110010111111011101",
    "111100101111000000110111",
    "111100101011101110000110",
    "111100101001001001101100",
    "111100100111010110001010",
    "111100100110010101111000",
    "111100100110001011001001",
    "111100100110111000001011",
    "111100101000011111000011",
    "111100101011000001101111",
    "111100101110100010000011",
    "111100110011000001101101",
    "111100111000100010001110",
    "111100111111000101000000",
    "111101000110101011010000",
    "111101001111010110000010",
    "111101011001000110001101",
    "111101100011111100011101",
    "111101101111111001010010",
    "111101111100111100111111",
    "111110001011000111101001",
    "111110011010011001001011",
    "111110101010110001010000",
    "111110111100001111010110",
    "111111001110110010101110",
    "111111100010011010011011",
    "111111110111000101010011",
    "000000001100110001111110",
    "000000100011011110110101",
    "000000111011001010000101",
    "000001010011110001101110",
    "000001101101010011100010",
    "000010000111101101000101",
    "000010100010111011110000",
    "000010111110111100110000",
    "000011011011101101000100",
    "000011111001001001100010",
    "000100010111001110110011",
    "000100110101111001010111",
    "000101010101000101100010",
    "000101110100101111100001",
    "000110010100110011010110",
    "000110110101001100111110",
    "000111010101111000001010",
    "000111110110110000101001",
    "001000010111110010000001",
    "001000111000110111110101",
    "001001011001111101100001",
    "001001111010111110100000",
    "001010011011110110001001",
    "001010111100011111110001",
    "001011011100110110101101",
    "001011111100110110010001",
    "001100011100011001110011",
    "001100111011011100101010",
    "001101011001111010001110",
    "001101110111101101111101",
    "001110010100110011010111",
    "001110110001000110000101",
    "001111001100100001110001",
    "001111100111000010001111",
    "010000000000100011011011",
    "010000011001000001010111",
    "010000110000011000010010",
    "010001000110100100100001",
    "010001011011100010100111",
    "010001101111001111010010",
    "010010000001100111011001",
    "010010010010101000000101",
    "010010100010001110100111",
    "010010110000011000100010",
    "010010111101000011100110",
    "010011001000001101110001",
    "010011010001110101010000",
    "010011011001111000100011",
    "010011100000010110010101",
    "010011100101001101100101",
    "010011101000011101100001",
    "010011101010000101101000");


signal sample : boolean := false;
signal sampled : boolean := false;

signal I_asynch, Q_asynch : signed (23 downto 0);

signal filtk : signed(23 downto 0);
signal prod : signed (47 downto 0);
signal mac_I : signed (65 downto 0);
signal mac_Q : signed (65 downto 0);
signal sample_data : signed(23 downto 0);
	
signal read_pointer_I, read_pointer_Q : integer range 0 to 257;
signal clk_out_next : boolean := false;

signal inbuffer : std_logic_vector(23 downto 0);
	
begin

sample_ff : process(clk_sample, sampled)
	begin
		if sampled = true then
			sample <= false;
		elsif clk_sample'event and clk_sample = '1' then
			inbuffer <= data_in;
			sample <= true;
		end if;
	end process;
	
I_asynch <= Ia(read_pointer_I);
Q_asynch <= Qa(read_pointer_Q);
			
downconversion : process (clk_in)
	variable n : integer range -1 to 500;
	variable ns : integer range 0 to 2;
	variable nn : integer range 0 to 247;
	variable m : integer range 0 to 31 := 0;
	variable p : integer range 0 to 800;
	variable write_pointer, write_pointer_last : integer range 0 to 257 := 0;
	
	begin	
		if clk_in'event and clk_in = '1' then		
			if clk_out_next = true then
				clk_out <= '1';
			else
				clk_out <= '0';
			end if;

			if sample = true then
				sampled <= true;			
			elsif sampled = true then
				sampled <= false;
				if m = 0 or m = 4 or m = 8 or m = 12 or m = 16 or m = 20 or m = 24 or m = 28 then
					Ia(write_pointer) <= signed(inbuffer);  				-- 1
					--Qa(write_pointer) <= to_signed(0,24); 		-- 0
					m := m + 1;
				elsif m = 1 or m = 5 or m = 9 or m = 13 or m = 17 or m = 21 or m = 25 or m = 29 then
					--Ia(write_pointer) <= to_signed(0,24);		-- 0
					Qa(write_pointer) <= signed(inbuffer);			-- 1
					m := m + 1;
					clk_out_next <= false;
				elsif m = 2 or m = 6 or m = 10 or m = 14 or m = 18 or m = 22 or m = 26 or m = 30 then
					Ia(write_pointer) <= signed(not inbuffer) + 1; -- -1
					--Qa(write_pointer) <= to_signed(0,24); 	 -- 0
					m := m + 1;
				elsif m = 3 or m = 7 or m = 11 or m = 15 or m = 19 or m = 23 or m = 27 or m = 31 then
					--Ia(write_pointer) <= to_signed(0,24);		-- 0
					Qa(write_pointer) <= signed(not inbuffer) + 1; -- -1

					if m = 31 then  -- clock out and start filter
						clk_out_next <= true;
						m := 0;    -- written samples
						n := -1;	  -- filter multiplication steps	
						ns := 2;	  
						prod <= to_signed(0,48);
						mac_I <= to_signed(0,66);
						mac_Q <= to_signed(0,66);	
						
						p := write_pointer_last;
						if p > 257 then
							read_pointer_I <= p - 258;
							read_pointer_Q <= p - 258;
						else
							read_pointer_I <= p;
							read_pointer_Q <= p;
						end if;
					else
						m := m + 1;
					end if;
					
				end if;
				
				if m = 0 or m = 2 or m = 4 or m = 6 or m = 8 or m = 10 or m = 12 or m = 14 or m = 16 or m = 18 or m = 20
							or m = 22 or m = 24 or m = 26 or m = 28 or m = 30 then	--- these are new m's		
					write_pointer_last := write_pointer;
					if write_pointer = 0 then
						write_pointer := 257;
					else
						write_pointer := write_pointer - 1;
					end if;
				end if;	
			end if;
			
			if not (m = 0 and sampled = true) then
				if n > -1 and n < 497 then
					if ns = 0 then  -- filtk and sample now for Q - compute prod for Q, prod now is for I
						sample_data <= I_asynch;
						mac_I <= mac_I + prod;
						p := read_pointer_Q + 1;
						if p > 257 then
								read_pointer_Q <= p - 258;
						else
							read_pointer_Q <= p;
						end if;
						ns := 1;
					elsif ns = 1 then
						sample_data <= Q_asynch;
						mac_Q <= mac_Q + prod;
						p := read_pointer_I + 1;
						if p > 257 then
							read_pointer_I <= p - 258;
						else
							read_pointer_I <= p;
						end if;
						ns := 0;
					end if;
					prod <= sample_data*filtk;
				end if;
				
				if n = -2 then
					n := -1;
				elsif n = -1 then
					filtk <= filtkoeff(0);
					sample_data <= Q_asynch;
					n := 0;
					ns := 0;  -- start with multiplication of Q
				elsif n < 495 then
					if n < 247 then
						nn := n + 1;   -- nn = 0 to 247
					else 
						nn := 494 - n; -- nn = 247 to 0, symmetric filter, only half of the taps need to be stored
					end if;
					filtk <= filtkoeff(nn);
					n := n + 1;
				elsif n = 495 or n = 496 then -- n = 495, final I mult and Q mac, n = 496 final Q mac
					n := n + 1;
				elsif n = 497 then
					if rx_att = "11" then
						Data_out_I <= std_logic_vector(mac_I + to_signed(268435456,60))(52 downto 29);  
						Data_out_Q <= std_logic_vector(mac_Q + to_signed(268435456,60))(52 downto 29);
					elsif rx_att = "10" then
						Data_out_I <= std_logic_vector(mac_I + to_signed(134217728,60))(51 downto 28); 
						Data_out_Q <= std_logic_vector(mac_Q + to_signed(134217728,60))(51 downto 28);
					elsif rx_att = "01" then
						Data_out_I <= std_logic_vector(mac_I + to_signed(67108864,60))(50 downto 27);  
						Data_out_Q <= std_logic_vector(mac_Q + to_signed(67108864,60))(50 downto 27);
					else
						Data_out_I <= std_logic_vector(mac_I + to_signed(33554432,60))(49 downto 26);  
						Data_out_Q <= std_logic_vector(mac_Q + to_signed(33554432,60))(49 downto 26);
					end if;	
					n := 498; -- to stop
				end if;
			end if;
		end if;
	end process;

end down_dec_arch;



library ieee;
use ieee.std_logic_1164.ALL;
use ieee.std_logic_unsigned.ALL;
use ieee.numeric_std.ALL;

entity down_dec_old is
	port (Data_in : in std_logic_vector(23 downto 0);
			Data_out_I : out std_logic_vector(23 downto 0);
			Data_out_Q : out std_logic_vector(23 downto 0);
			clk_in : in std_logic; -- 40 MHz
			clk_sample : in std_logic; -- 40 / 32 MHz
			rx_att : in std_logic_vector(1 downto 0);
			clk_out : out std_logic
			);
end down_dec_old;

architecture down_dec_arch of down_dec_old is

--signal Data_in_trunk : signed (17 downto 0);
-- signal Ia : signed (8 downto 0);
-- signal Qa : signed (8 downto 0);
--signal mac_I_sig : signed (23 downto 0);
--signal mac_Q_sig : signed (23 downto 0);
	
type longbuffer is array (200 downto 0) of signed (23 downto 0);
type filt_type is array (159 downto 0) of signed (23 downto 0);

signal Ia : longbuffer;
signal Qa : longbuffer;

constant filtkoeff : filt_type :=

-- Scilab:
-->[v,a,f] = wfir ('lp', 160, [1/120 0], 'hn', 0);
-->round(v*2^28)

	("000000000000000000000000",
    "111111111111111010100010",
    "111111111111101010101011",
    "111111111111010001011011",
    "111111111110110000000011",
    "111111111110001000000000",
    "111111111101011010111111",
    "111111111100101010111011",
    "111111111011111001111100",
    "111111111011001010011001",
    "111111111010011110110010",
    "111111111001111001110110",
    "111111111001011110011010",
    "111111111001001111011111",
    "111111111001010000001110",
    "111111111001100011110101",
    "111111111010001101101010",
    "111111111011010001000101",
    "111111111100110001011111",
    "111111111110110010010110",
    "000000000001010111000011",
    "000000000100100010111111",
    "000000001000011001011111",
    "000000001100111101110000",
    "000000010010010010111011",
    "000000011000011011111110",
    "000000011111011011101011",
    "000000100111010100101011",
    "000000110000001001010110",
    "000000111001111011110110",
    "000001000100101110000110",
    "000001010000100001101100",
    "000001011101010111111100",
    "000001101011010001110101",
    "000001111010010000000010",
    "000010001010010010110101",
    "000010011011011010001011",
    "000010101101100101101001",
    "000011000000110100011001",
    "000011010101000101010000",
    "000011101010010110100111",
    "000100000000100110011111",
    "000100010111110010100000",
    "000100101111110111111001",
    "000101001000110011100001",
    "000101100010100001111000",
    "000101111100111111000100",
    "000110011000000110111000",
    "000110110011110100110000",
    "000111010000000011110100",
    "000111101100101110111010",
    "001000001001110000100110",
    "001000100111000011001100",
    "001001000100100000110011",
    "001001100010000011010100",
    "001001111111100100011111",
    "001010011100111101111011",
    "001010111010001001000111",
    "001011010110111111011111",
    "001011110011011010011101",
    "001100001111010011011001",
    "001100101010100011110000",
    "001101000101000101000000",
    "001101011110110000110000",
    "001101110111100000101101",
    "001110001111001110110010",
    "001110100101110101000011",
    "001110111011001101110110",
    "001111001111010011110000",
    "001111100010000001101010",
    "001111110011010010110001",
    "010000000011000010100111",
    "010000010001001101001001",
    "010000011101101110101001",
    "010000101000100011110111",
    "010000110001101001111101",
    "010000111000111110100010",
    "010000111110011111101010",
    "010001000010001011111001",
    "010001000100000010010001",
    "010001000100000010010001",
    "010001000010001011111001",
    "010000111110011111101010",
    "010000111000111110100010",
    "010000110001101001111101",
    "010000101000100011110111",
    "010000011101101110101001",
    "010000010001001101001001",
    "010000000011000010100111",
    "001111110011010010110001",
    "001111100010000001101010",
    "001111001111010011110000",
    "001110111011001101110110",
    "001110100101110101000011",
    "001110001111001110110010",
    "001101110111100000101101",
    "001101011110110000110000",
    "001101000101000101000000",
    "001100101010100011110000",
    "001100001111010011011001",
    "001011110011011010011101",
    "001011010110111111011111",
    "001010111010001001000111",
    "001010011100111101111011",
    "001001111111100100011111",
    "001001100010000011010100",
    "001001000100100000110011",
    "001000100111000011001100",
    "001000001001110000100110",
    "000111101100101110111010",
    "000111010000000011110100",
    "000110110011110100110000",
    "000110011000000110111000",
    "000101111100111111000100",
    "000101100010100001111000",
    "000101001000110011100001",
    "000100101111110111111001",
    "000100010111110010100000",
    "000100000000100110011111",
    "000011101010010110100111",
    "000011010101000101010000",
    "000011000000110100011001",
    "000010101101100101101001",
    "000010011011011010001011",
    "000010001010010010110101",
    "000001111010010000000010",
    "000001101011010001110101",
    "000001011101010111111100",
    "000001010000100001101100",
    "000001000100101110000110",
    "000000111001111011110110",
    "000000110000001001010110",
    "000000100111010100101011",
    "000000011111011011101011",
    "000000011000011011111110",
    "000000010010010010111011",
    "000000001100111101110000",
    "000000001000011001011111",
    "000000000100100010111111",
    "000000000001010111000011",
    "111111111110110010010110",
    "111111111100110001011111",
    "111111111011010001000101",
    "111111111010001101101010",
    "111111111001100011110101",
    "111111111001010000001110",
    "111111111001001111011111",
    "111111111001011110011010",
    "111111111001111001110110",
    "111111111010011110110010",
    "111111111011001010011001",
    "111111111011111001111100",
    "111111111100101010111011",
    "111111111101011010111111",
    "111111111110001000000000",
    "111111111110110000000011",
    "111111111111010001011011",
    "111111111111101010101011",
    "111111111111111010100010",
    "000000000000000000000000");

--attribute ramstyle : string;
--attribute ramstyle of filtkoeff : constant is "M4K";

signal sample : boolean := false;
signal ack : boolean := false;

signal I_asynch,Q_asynch, I_synch, Q_synch : signed (23 downto 0);

signal mac_I : signed (60 downto 0);
signal mac_Q : signed (60 downto 0);

signal write_pointer, write_pointer_last : integer range 0 to 255 := 200;
signal read_pointer : integer range 0 to 255;
signal clk_out_next : boolean := false;
	
begin

downconversion : process (clk_in)
	variable ns : integer range 0 to 3 := 0;	
	begin	
		if clk_in'event and clk_in = '1' then		
			if clk_out_next = true then
				clk_out <= '1';
			else
				clk_out <= '0';
			end if;

			if sample = true then
				ack <= true;
				if ns = 0 then
					Ia(write_pointer) <= signed(Data_in);  				-- 1
					Qa(write_pointer) <= to_signed(0,24); 		-- 0
					ns := 1;
				elsif ns = 1 then
					Ia(write_pointer) <= to_signed(0,24);		-- 0
					Qa(write_pointer) <= signed(Data_in);			-- 1
					ns := 2;
				elsif ns = 2 then
					Ia(write_pointer) <= (not signed(Data_in)) + 1; -- -1
					Qa(write_pointer) <= to_signed(0,24); 	 -- 0
					ns := 3;
				elsif ns = 3 then
					Ia(write_pointer) <= to_signed(0,24);		-- 0
					Qa(write_pointer) <= (not signed(Data_in)) + 1; -- -1
					ns := 0;
				end if;		
				write_pointer_last <= write_pointer;
			else
				ack <= false;
			end if;
			I_asynch <= Ia(read_pointer);
			Q_asynch <= Qa(read_pointer);
			I_synch <= I_asynch;
			Q_synch <= Q_asynch;
		end if;
	end process;
	
filter : process (clk_in)
	variable prod_I : signed (47 downto 0);
	variable prod_Q : signed (47 downto 0);
	variable n, nn : integer range 0 to 160 := 0;
	variable m : integer range 0 to 31 := 0;
	variable filter_start_pointer : integer range 0 to 200 := 100;
	variable p : integer range 0 to 511;

	begin	
		if clk_in'event and clk_in = '0' then
			if ack = true then	
				if write_pointer = 0 or write_pointer > 200 then
					write_pointer <= 200;
				else
					write_pointer <= write_pointer - 1;
				end if;		
				if m = 31 then
					filter_start_pointer := write_pointer_last;
					m := 0;
					n := 0;			
				else
					m := m + 1;
				end if;
			end if;

			p := filter_start_pointer + n;
			if p > 200 then
				read_pointer <= p - 201;
			else
				read_pointer <= p;
			end if;
			
			if n < 160 then
				if n = 1 then
					nn := 159;
				elsif n = 0 then
					nn := 158;
				else
					nn := n - 2;
				end if;
				
            prod_I := I_synch*filtkoeff(nn);  -- Ia(32*m)
				prod_Q := Q_synch*filtkoeff(nn);
				
				if nn = 0 then
					if rx_att = "11" then
						Data_out_I <= std_logic_vector(mac_I + to_signed(268435456,60))(52 downto 29);  
						Data_out_Q <= std_logic_vector(mac_Q + to_signed(268435456,60))(52 downto 29);
					elsif rx_att = "10" then
						Data_out_I <= std_logic_vector(mac_I + to_signed(134217728,60))(51 downto 28); 
						Data_out_Q <= std_logic_vector(mac_Q + to_signed(134217728,60))(51 downto 28);
					elsif rx_att = "01" then
						Data_out_I <= std_logic_vector(mac_I + to_signed(67108864,60))(50 downto 27);  
						Data_out_Q <= std_logic_vector(mac_Q + to_signed(67108864,60))(50 downto 27);
					else
						Data_out_I <= std_logic_vector(mac_I + to_signed(33554432,60))(49 downto 26);  
						Data_out_Q <= std_logic_vector(mac_Q + to_signed(33554432,60))(49 downto 26);
					end if;
					mac_I <= to_signed(0,61) + prod_I;
					mac_Q <= to_signed(0,61) + prod_Q;
				else
					mac_I <= mac_I + prod_I;
					mac_Q <= mac_Q + prod_Q;
				end if;
				
				if nn = 2 then
					clk_out_next <= true;
				else
					clk_out_next <= false;
				end if;

            n := n + 1;
         end if;
			
		end if;
	end process;
	
	sample_ff : process(clk_sample,ack)
	begin
		if ack = true then
			sample <= false;
		elsif clk_sample'event and clk_sample = '1' then
			sample <= true;
		end if;
	end process;
	
end down_dec_arch;